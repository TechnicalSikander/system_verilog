`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: IIT JAMMU
// Engineer: Mohammad Sikander Sheikh
// 
// Create Date: 01.09.2025 23:28:24
// Design Name: 
// Module Name: two_port_ram
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: it is not infer the BRAM it infer the LUT
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module two_port_ram
#(parameter A_WIDTH = 3 , D_WIDTH = 8)
(
input logic clk, we,
input logic [A_WIDTH -1 :0] r_add,
input logic [A_WIDTH -1 :0] w_add,
input logic [D_WIDTH -1 :0] w_data,
output logic [D_WIDTH -1 : 0] r_data
    );

logic [D_WIDTH - 1 : 0 ] mem[0:2**A_WIDTH -1];
//write
always_ff@(posedge clk)
begin
 if(we)
   mem[w_add] <= w_data;
 end
 assign r_data = mem[r_add];

endmodule
